isrc 1 0 0.0 0.0 1.0e-9 0.5e-3 2.0e-9 0.25e-3 3.0e-9 0.0 4.0e-9 0.0
res 1 2 100.0
cap 1 0 1.0e-12
cap 2 0 3.0e-12
