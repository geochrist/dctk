isrc 1 0 0.0 0.0 1.0e-9 0.5e-3 2.0e-9 0.25e-3 3.0e-9 0.0 4.0e-9 0.0
res 1 2 100.0
cap 1 0 1.0e-12
cap 2 0 3.0e-12
res 1 3 150.0
cap 3 0 1.75e-12
res 3 4 125.0
cap 4 0 2.5e-12
res 4 5 75.0
cap 5 0 3.75e-12
